       I              �iW�
�@                     q       e        Icarus Verilog                                                                                                                  Tue Apr 15 14:40:52 2025
                                                                                                             �              �      ���
ex^���`��Q@m  ��?eZ ���������!x^c�   ���x^c`c��p�B �L]  �x^c`� ���l��Т��  Q A5x^c�p��R��  44�  Q�  �  ��   n�
   ��x^c�� A.0�gY 
�O   j0 �x^c�  ظ��
�����*�턕�T�04-f&�h H)�p1� �b��,�X�aQ�2A�< U`��lb �&b}�H�OF���������������������OnKH����@U �G�?0x^c�  �� �׊�X �)�x^��!� PJ*J�@LLLL� o��N�I��M���A~�����W:?�5Ucɐ���P-c���	]���E��)�r\� m���ٸ_��y�����&��M>����J�Nix^c�p��pR��h�z��ox^c`s��P2����B �F�x^c```bd�@,,�`R ���"C|Td0� I �	?^�x^�ʱ�0C��
R��d��2#0#0�B��
qe=X�O|����r�*C7��(�ҫuw6�r�C��2|���M��x �vdάx^c�  ظ��
00m`hZ�,� \,,��Y� â&et�Q.��� t�v7�x^퓱�0?ȅ)RPPPP0��c)v�I¿B�(�N�|'w���x�Ĝ� ȎH���^t31C�]� ��dcw7��ڞ���򺃝$�@mO   �x^c`�B-0��) �	�x^c` n(��
X�Jր�j����` "x�\�,��`���H��`���I��q Y2�:�:@J8@:�&��U7�n�S` Umf xxxxxxxx X�   �  ����������  j� �@|�  n� �@|��x^c`(�``�`Q`�`1`�`q`�`	`�`I`�`)`�`i`�`��2�e�
�,;X��`��r����,?XXF���@? ��o   �� �0�@�P�`�p��   n��V�+��
���� �x^c�  ��@����A��2�bÙ�  %�c�x^cp�R��ВP�P�Аq	t�  ���kx^c�����" ��!��  |��ox^c� >�"4h��6  ��"��x^c� �	  �� ٷ�px^c� � 	 �4�  ��x^c�  ���,�0 ��00H0��< 1	�O� ���H�G%F%K  �S2��x^c�  ���000�K��R����,���`�sY\@� �,�`�DΈf���Q����Q��I֎�g _"�rx^c� � �
" ��� T� ��x^c�  �X8�� ��@B$&$@b2"@B$� BD�J�J�"&4 ��"{�x^c�  ���20p 	F0�$�@�� �p� q�< BD�� 	9K	�N�N.�1*;*;dd�\ ��A=�x^c````ab@�D��	 !bI� � SsA�(��\ ��~�x^c�  ��� 	 �`a`0��@#�����$X@, Y	�,H�!H�UۨĨa	D�b �����x^c�@�@ a������,F�1����,f�fa`�Y��R,�!�Q,�"�X�IC��Ih� ��,����y�ZȈ��Qm�2��0dF�aȌjÐ��6E%C1�C1 Mjȥx^햱� E��&�v.`\���U�C<��1�Cl�����BG1
��=��ku�{�*G�����B��RDy `#Jpމ��me�RX-�;�dC�:�(�,7[�Y,��7�D%BT����=*Q�7���O(1�6����x^c4��
(`G@�X�Up0��0a�����!�������� �!��P�� ���AC(���(�K�0X^��a1�$PN;G��j�6�m�j#��,�"�  Z@n�x^c�  ���� �0 ��a�``�p�� HL.�1
�X,��G%F%K  ��#� � �(  �(�5x^c�ĨP�D 7��4x^cq2�2p"	 (�` 5x^cSR�bR  1%� " px^c�� ..�6@�AC �)!آx^c����bHp�x � � ��  R�&��x^c� ����������?,�D�����$��`��`55`Y���	 �	�����M(����7  g1䭬x^c�  ��
 	�!$�\.L�Q.��� T�Q�x^c�  ��� 	 �`a`0��@#\�$�% ����2�dA����F%F%K # �W!	Qx^c��P�0�%��  �U�;x^c��P�0�I�Y$@� J��6x^c��RRH��")  2���x^c��� �U Ѵ�A�A��A�� ����A]l�K#.0
 �W_�x^c�  �V	 	V������� �
wd� ;Qy�x^c���X9�00000-��``�`��Y����%�!6ʥ��� �_{K�x^c�  ��
 	�!$���� ����҈� -�v�x^c���V	00p� 	6����� �XDP�#��  ��x��x^c�  ��� 	 fd�L���2��1Ȁ$@JJ$Fņ�(j���Ox^c���P�RR0� �iάx^c�  ����
00m`hZ�,� \,,��Y� â&et�Q.��� { v;�x^c` &F ! $X@���  ���2 10D�r��U �y>�x^c``S`q`I`a`A�X`���D���C��-�  Ie]�      )%� 	)/�-u�15� �}� �1_K�g!	m� �7;� ac� 1=�=;� �9� �_]� ����� '�~%%�~5� �� �11-� � � � � � /� �_� � �       �x�c��`� J��      �             �       Y       e       ex�M�1
�0���;���?Y�Yr2HB`!YMVv�7<��jD8��\����k|�a�m~��]      W      x�      
}TYo�@^'�@�<!�P�8����C�U%GU)A+�ɪ>���I�{�2���ni#�3�������H7<^~��"	S�/�pr9r�9��~�C*�����"�������B�dvE,��\��,F��ɀ�ď��	�|����#�Q:�C��	��[:��7�����{`a9�<�� �w��A<���'���t"Z��4� K�Z���֦����=$	�ɅG�<�*o���_Sf��`�
�f5/�G���B��%!�e�Tp�k`>�̴<�8��d�K��)�3A#�@��蓒W����@tJgW4#��'��*Э�@;d�D�����k�^��"��a��8��7D�xE��~�q]��ϼ-ϴY�k���^��<�����{�~Ӈ�/Q��S�d����� ��}R�.�%�Q���zL�Ң �_�j�Q� ��|)li�4��Cgï�KW�ϊT���e��P�,XCU�D�B���k�'X�#�%0���&��� �Ju��Cs�j��T�r�J���n����zR�W
$����ƣ�r#�F�aCp��u�r�vQ1���`��j�X�H������ڸ|�Sl�y �kʒ�!z�.�=��Ni�Ȩ�W������8ژ+������N�q2�����Q��Z�eH@�Z�HZ����k�����@�SZ=�W��l|�6���8�#ߤ�/��Ϙ�3�`� �%�&�wr�RR���l.�(������i8k�m�k��x�&d56a���q�:�vp�@�`J�,b�F�6Y���w��݌W���{���W�x  