       I            .��iW�
�@                     �       �       �Icarus Verilog                                                                                                                  Fri Apr 18 20:54:46 2025
                                                                                                             �            .��      �	��x^���`��Q0
F�� ��F�Z !x^c�   �� ���������Sx^��1  ���K��^�         �BȁЙ  R   /xxxx  �  �    �   �
   ���@���P�(���J��  � Ta   7xxxx+x^c` &F �[A   ��1 �      �
     -xxxxxxxxxxxxxxxx      �
             /xxxxxxxxxxxx     /xxxxxxxxxxxxxxxxxxxxxxxx  Pa$x^c` }(��
 �-  �z�������� ���������  ��  P> �@��   �� �0�@�P�`�p�� xxxxxP@ �@���x^c� 6� 	� ����|�,,,Xf�,`Y���e��,Xn�<`y���Ǩ��� �	�0 xxxxxxxx��x^��1  0�rW9��Z�c�!Yrz��V_۶m۶m۶m۶m۶m۶m۶m۶m۶m۶m���[N��x^��1  0�rW9��X�c�!Yrz��V_۶m۶m۶m۶m۶m۶m۶m۶m۶m۶m��giL�   �     xxxx xxxxx        xxxxxxxxxxxxxxxx 00000000xxxxxxxx xxxxxxx xxx xxxxxxxxxxxx"x^c�  Kz!x^c���  ���!x^c�� �z�            * 00xx0       xxxxxxxxP�Wx^c�  .02 A�d�L`�L��IV0�&��$ �k�%� s	g	7		}s)os	1}Cg#Y=}g%?=_7'�]g�C}���Ag�~}Y�~�~�~�~}�~�~}C�~}Sg}%�~%}�~}�}}����~��~}       �x���  ����c��1�                    �(�m      Sq       .      )�       i       �       �x�MMA�0
�dz�q������.]�� Q� 2�$�rH]j��g'#ɜ�4G��JP�IЮG�<�pa��ԟ�ӎR��z���      �      ��      
�W�n7�JZ��6�C�
衧�^������ue90`��P���W�k�}���y-C���%W��̷����}G�����2�sVHq���Ip)x|)#*������#O��~o	�TF����t���sZ�w'��iyx19z������������'qv��r!i������ ����o���%�6~���X���2Kh�@ ���B�4t6��A��njě0KZ1�V+��L�Mp���!��y�Zo6���.~�t��IY0�jq�|��v�����%F��A���,�k�@��]5�5M�s#��2��a���A�$�.
�iθ�J�
�r�!�F>=�q>�Ո��o��u�e�έ�5�_Ȓ�JI�)� �G? 8��Xp������a��`�?%N�zcq�C�~���aQ�mh��!(���28�BB!��E�x{�n1�P�<�r�,~I4��Z���KnN��k�j���w�uƝ
�_�؛���G�H�nj�=Ŧ��]x��i��{��%TV|-��e�e}�D�Ԁ��)�l#������@�Ǔ�4.�Ғ�>�k?"�>�Iߌ���������"��@��-�$R� ���f�$��y�W}f�C׬fʢơ��>�Yxn|mKk����?���O.�:�\���i��m�k�f�9��; ��[�:���Qì��ȹ�-�Mp�r�)���Rܡ��d��3��䣻���[T�H�iU���Vtnemq���Zfz؀�s�t�IV��M镎�ᆭ��N'Ú
P-��UL�:2�S#� CM�7,�%���)@gʪeS��\���v�	-�'�ߌ��ҝ��
*o�.��MG���Acz�����b�; ��G�<�G_8�I82��
^���B��G�{�ãS5hm����jL��R��n�J/v��=�ڤ�-�n�vZ+��&�&�r��D�\� 6:z2r��"^�gm��
4���������
d#Naɉ~,�"�//~Ġ�`�N��:�Y@�?�U#�#X��~m��ވl�Cǋ3��[��?�x֯��>����k�}h�6�:S�M��(��=�~��z 5�r|>�`��>�]�qRt�Ƿ����^ ������������X�����^����YZM�6ݢ���G��8�o=5It^]��=x��Ph�p�  