       I              ^iW�
�@                                    Icarus Verilog                                                                                                                  Fri Dec 06 01:39:57 2024
                                                                                                             [              ^      15x^��   ��Z �  �  ��x^c`c��p� ��� xxxxxxxx     �  ����������  � �@|�  � �@|��x^c`��``�`Q`�`1`�`q`�`	`�`I`�`)`�`i`�`��2�e�
�,;X��`��r����,?XXF���@? ��   �� �0�@�P�`�p��   'w		{}� �7       x�c��`� G�_      $             $       )                          ��      
u��J�0�/]#~�<@�	¾)>��"�r�i&e���"���f.���������e�Y�,�z�?lG�4v���-�`J��끐��/Hr�<�;x~XX<(�Du�٘T�}�D�i�1֚�|}��y��P:�����'t���pP�A��������K[�T���S�1KB�Ʒmpê!wOBc�\��ش�=��^Ǫ�#�#Mv��c��������wd��zd�n�q�]���OO���� �">_�  