       I             A'�iW�
�@                                   �Icarus Verilog                                                                                                                  Fri Apr 18 19:42:35 2025
                                                                                                             �             A'�      [x^���  ��*�Z  ��   ���@���P�(���J���x^c`c��pR �(� ��������  � �z�������� ���������  ��  �> �@���   �� �0�@�P�`�p���  xxxxx�@ �@����x^c� 6�F	� ����|�,,,Xf�,`Y���e��,Xn�<`y���Ǩ��� ��a xxxxxxxx��Wx^c�  ����H0�I&0�&Y�$+�d��`� ���7)%}?=#=/�       x�c�P��p��Q8
7 �lG�      �             W       )                           ��      
u��j�0��1�1�h�`l��s�`�]�a�e�Y�R�w�,'����e��'i���cc�o[�ˌ}��m3ך�r��T�?_ H������r �EWe��&�����'!a���%�>������?�F]y�
b�1�{�b=�T��b��J3�rMM�"Ɨ�N�Jsva�SWU����KbA��=)G�l��1G�u�A���ɶI��B4�.�JS�y��6{s��1�g.������u�����@����$�_����  